//第２回計算機システム設計論演習問題(1-2)

module test(a,b);
	output b;
	input a;
	assign b = a;
endmodule